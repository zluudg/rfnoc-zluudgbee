----------------------------------------------------------------------------------------------------
-- Project: IT245X Degree Project in Microelectronics
-- Developer: Leon Fernandez
-- Component: decimator ("Keep one in N"-style decimator)
-- Description: Will let through every N:th packet, determined by
-- one of the input. Additionally, it has an input to adjust the offset.
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.zluudg_constants.all;

entity zluudg_decimator is
    port ( aclk               : in std_logic;
           areset             : in std_logic;
           shift              : in std_logic_vector(1 downto 0);
           sr_decim_rate      : in std_logic_vector(C_SETREGW - 1 downto 0);
           s_iqsample_tready  : out std_logic;
           s_iqsample_tvalid  : in std_logic;
           s_iqsample_tlast   : in std_logic;
           s_iqsample_tdata	  : in std_logic_vector(C_IQSAMPLEW - 1 downto 0);
           m_tready           : in std_logic;
           m_tvalid           : out std_logic;
           m_sym_tdata        : out std_logic_vector(C_IQSAMPLEW - 1 downto 0);
           m_oldsym_tdata     : out std_logic_vector(C_IQSAMPLEW - 1 downto 0));
end zluudg_decimator;

architecture Behavioral of zluudg_decimator is

    -- Delay data signal two cycles to match the delay in
    -- calculating the error signal. This way, the value of
    -- the error signal corresponds to the current value
    -- being output
    signal tdata_d : std_logic_vector(C_IQSAMPLEW - 1 downto 0) := (others => '0');

    -- Delay blip from "en_decim" for use as output tvalid. The delay is needed
    -- since the output is delayed by two cycles.
    signal tvalid_d : std_logic := '0';

    -- The previous decimated symbol that we let through
    signal prev_symbol : std_logic_vector(C_IQSAMPLEW - 1 downto 0) := (others => '0');

    -- Treat both input tready signals as one signal
    signal m_axis_tready : std_logic;

    -- Counter that counts upwards and wraps around whenever a decimation is performed
    signal counter : unsigned(C_DECIM_COUNTERW - 1 downto 0) := (others => '0');

    -- Counter that takes into account whether we are shifting this cycle or not
    signal decim_counter : unsigned(C_DECIM_COUNTERW - 1 downto 0) := (others => '0');

    -- Typecast version of the input shift signal for easy addition
    signal shift_arith : unsigned(1 downto 0);

    -- Enable signal for the output register
    signal en_decim : std_logic := '0';

begin

    -- This block is always ready if the succeeding blocks are ready and it is not resetting.
    s_iqsample_tready <= m_tready and (not areset);

    -- The registered input drives the output and "m_tvalid" is used to pass a subset
    -- of the input samples to the next block.
    m_sym_tdata <= tdata_d;

    -- The prev_symbol register stores the previous decimated sample that was flagged with
    -- "m_tvalid". The conjugate of that previous sample is then output on the
    -- "oldsym" AXIS master interface.
    m_oldsym_tdata(C_IQSAMPLEW - 1 downto C_SAMPLEW) <=
        std_logic_vector(-signed(prev_symbol(C_IQSAMPLEW - 1 downto C_SAMPLEW)));
    m_oldsym_tdata(C_SAMPLEW - 1 downto 0) <= prev_symbol(C_SAMPLEW - 1 downto 0);

    -- The counter used for decimation is the regular counter + the shift
    shift_arith <= unsigned(shift);
    decim_counter <= counter + shift_arith;

    -- The "m_tvalid" flags generated by the decimation counter
    m_tvalid <= tvalid_d;

    -- Feed through all data, use "valid" signal to mark desired symbols.
    P_TDATA_DLY: process (aclk)
    begin
        if rising_edge(aclk) then
            if (areset = '1') then
                tdata_d <= (others => '0');
            else
                if (s_iqsample_tvalid = '1' and en_decim = '1') then
                    tdata_d <= s_iqsample_tdata;
                end if;
            end if;
        end if;
    end process P_TDATA_DLY;


    -- A process that uses the "m_tvalid" flag generated by the decimation
    -- counter to store the previous valid symbol in a register that drives
    -- the "oldsym"-output.
    P_OLDSYM: process (aclk)
    begin
        if rising_edge(aclk) then
            if (areset = '1') then
                prev_symbol <= (others => '0');
            else
                if (tvalid_d = '1') then
                    prev_symbol <= tdata_d;
                end if;
            end if;
        end if;
    end process P_OLDSYM;
    
    -- A counter that asserts a signal every DECIMATION_RATE:th input.
    -- This signal drives the tvalid flags on the master/output interfaces.
    -- If the "shift" signal is asserted, this counter asserts a signal
    -- every "DECIMATION_RATE-1":th input until the "shift" signal is
    -- deasserted.
    P_DECIM_COUNTER: process (aclk)
    begin
        if rising_edge(aclk) then
            if (areset = '1') then
                counter <= (others => '0');
                en_decim <= '0';
            else
                if (s_iqsample_tvalid = '1') then
                    if (decim_counter = unsigned(sr_decim_rate)-1) then
                        en_decim <= '1';
                        counter <= counter + 1;
                    elsif (decim_counter = unsigned(sr_decim_rate)) then
                        en_decim <= '0';
                        counter <= (0=>'1', others => '0');
                    else
                        counter <= counter + 1;
                    end if;
                end if;
            end if;
        end if;
    end process P_DECIM_COUNTER;

    -- Process that delays the tvalid by one cycle to match the delay caused
    -- by the input register.
    P_TVALID_DLY: process (aclk)
    begin
        if rising_edge(aclk) then
            if (areset = '1') then
                tvalid_d <= '0';
            else
                tvalid_d <= en_decim and s_iqsample_tvalid;
            end if;
        end if;
    end process P_TVALID_DLY;

end Behavioral;